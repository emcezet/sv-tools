these are valid ids /* A block comment started,
we can use any keywords here like and or module
and the comment may be very very very very very
very very very very very very very very very very
very very very very very very very very very very
very very very very very very very very very very
very very very very very very very very very very
very very very very very very very very very very
very very very very very very very very very very
very very very very very very very very very very
long*/ again these are valid ids
/* Another block comment started,to check for
non greedy regexps expansion */
